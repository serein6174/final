`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/04/09 02:04:58
// Design Name: 
// Module Name: counter_1s
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module clk_2s(clk, clk_2s);
input wire clk;
output reg clk_2s;
reg [31:0] cnt;
always @ (posedge clk) begin
   
end
endmodule

