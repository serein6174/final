module digit(
    input [3:0] digit,  //����0-9
    input [3:0] row,     //�е�ַ0-15
    output reg [11:0] pixels //12λ�������ݣ������ң�
);
    always @(*) begin
        case({digit, row})
            //---------------- ���� 0 -----------------
            8'h00: pixels = 12'b000011110000;  
            8'h01: pixels = 12'b000111111000;
            8'h02: pixels = 12'b001111111100; 
            8'h03: pixels = 12'b011100011110; 
            8'h04: pixels = 12'b011000001110; 
            8'h05: pixels = 12'b111000001111;
            8'h06: pixels = 12'b111000000111; 
            8'h07: pixels = 12'b111000001111; 
            8'h08: pixels = 12'b011000001110; 
            8'h09: pixels = 12'b011100011110; 
            8'h0A: pixels = 12'b001111111100;
            8'h0B: pixels = 12'b000111111000; 
            8'h0C: pixels = 12'b000011110000;   
            8'h0D: pixels = 12'b000000000000;
            8'h0E: pixels = 12'b000000000000; 
            8'h0F: pixels = 12'b000000000000; 

            //---------------- ���� 1 -----------------
            8'h10: pixels = 12'b000000110000;   
            8'h11: pixels = 12'b000001110000;   
            8'h12: pixels = 12'b000011110000;  
            8'h13: pixels = 12'b000000110000;   
            8'h14: pixels = 12'b000000110000;  
            8'h15: pixels = 12'b000000110000;  
            8'h16: pixels = 12'b000000110000;    
            8'h17: pixels = 12'b000000110000;     
            8'h18: pixels = 12'b000000110000; 
            8'h19: pixels = 12'b000000110000;  
            8'h1A: pixels = 12'b000000110000;    
            8'h1B: pixels = 12'b000111111110; 
            8'h1C: pixels = 12'b000111111110;  
            8'h1D: pixels = 12'b000000000000;            
            8'h1E: pixels = 12'b000000000000; 
            8'h1F: pixels = 12'b000000000000; 

            //---------------- ���� 2 -----------------
            8'h20: pixels = 12'b000111111000; 
            8'h21: pixels = 12'b001111111100; 
            8'h22: pixels = 12'b011100011110; 
            8'h23: pixels = 12'b011000001110; 
            8'h24: pixels = 12'b000000001110; 
            8'h25: pixels = 12'b000000011100; 
            8'h26: pixels = 12'b000000111000;  
            8'h27: pixels = 12'b000001110000;     
            8'h28: pixels = 12'b000011100000;    
            8'h29: pixels = 12'b000111000000;     
            8'h2A: pixels = 12'b001111111110; 
            8'h2B: pixels = 12'b011111111110; 
            8'h2C: pixels = 12'b011111111110; 
            8'h2D: pixels = 12'b000000000000;             
            8'h2E: pixels = 12'b000000000000;            
            8'h2F: pixels = 12'b000000000000; 

            //---------------- ���� 3 -----------------
            8'h30: pixels = 12'b001111111000; 
            8'h31: pixels = 12'b011111111100; 
            8'h32: pixels = 12'b011000011100;
            8'h33: pixels = 12'b000000001110; 
            8'h34: pixels = 12'b000001111100;  
            8'h35: pixels = 12'b000001111100;   
            8'h36: pixels = 12'b000000001110; 
            8'h37: pixels = 12'b000000000110; 
            8'h38: pixels = 12'b000000000110; 
            8'h39: pixels = 12'b011000001110; 
            8'h3A: pixels = 12'b011111111100; 
            8'h3B: pixels = 12'b001111111000;
            8'h3C: pixels = 12'b000011100000;          
            8'h3D: pixels = 12'b000000000000;           
            8'h3E: pixels = 12'b000000000000;           
            8'h3F: pixels = 12'b000000000000; 

            //---------------- ���� 4 -----------------
            8'h40: pixels = 12'b000000011100;  
            8'h41: pixels = 12'b000000111100; 
            8'h42: pixels = 12'b000001111100; 
            8'h43: pixels = 12'b000011101100; 
            8'h44: pixels = 12'b000111001100; 
            8'h45: pixels = 12'b001110001100;  
            8'h46: pixels = 12'b011111111111; 
            8'h47: pixels = 12'b011111111111;
            8'h48: pixels = 12'b000000001100;
            8'h49: pixels = 12'b000000001100;  
            8'h4A: pixels = 12'b000000001100;  
            8'h4B: pixels = 12'b000000001100;  
            8'h4C: pixels = 12'b000000001100; 
            8'h4D: pixels = 12'b000000000000;          
            8'h4E: pixels = 12'b000000000000;            
            8'h4F: pixels = 12'b000000000000; 

            //---------------- ���� 5 -----------------
            8'h50: pixels = 12'b011111111110; 
            8'h51: pixels = 12'b011111111110; 
            8'h52: pixels = 12'b011000000000;         
            8'h53: pixels = 12'b011000000000;          
            8'h54: pixels = 12'b011111111000;     
            8'h55: pixels = 12'b011111111100;   
            8'h56: pixels = 12'b000000011110;         
            8'h57: pixels = 12'b000000001110;          
            8'h58: pixels = 12'b000000000110;           
            8'h59: pixels = 12'b000000001110;          
            8'h5A: pixels = 12'b011000011110;      
            8'h5B: pixels = 12'b011111111100;   
            8'h5C: pixels = 12'b001111111000;      
            8'h5D: pixels = 12'b000000000000;            
            8'h5E: pixels = 12'b000000000000;            
            8'h5F: pixels = 12'b000000000000; 

            //---------------- ���� 6 -----------------
            8'h60: pixels = 12'b000011111000;        
            8'h61: pixels = 12'b001111111100;    
            8'h62: pixels = 12'b011100001110;      
            8'h63: pixels = 12'b011000000110;        
            8'h64: pixels = 12'b011000000000;           
            8'h65: pixels = 12'b011011111000;      
            8'h66: pixels = 12'b011111111100;   
            8'h67: pixels = 12'b011110001110;     
            8'h68: pixels = 12'b011000000110;        
            8'h69: pixels = 12'b011000000110;        
            8'h6A: pixels = 12'b011100001110;      
            8'h6B: pixels = 12'b001111111100;    
            8'h6C: pixels = 12'b000011111000;        
            8'h6D: pixels = 12'b000000000000;          
            8'h6E: pixels = 12'b000000000000;         
            8'h6F: pixels = 12'b000000000000; 

            //---------------- ���� 7 -----------------
            8'h70: pixels = 12'b011111111110; 
            8'h71: pixels = 12'b011111111110; 
            8'h72: pixels = 12'b000000001110; 
            8'h73: pixels = 12'b000000011100;  
            8'h74: pixels = 12'b000000111000; 
            8'h75: pixels = 12'b000001110000;  
            8'h76: pixels = 12'b000011100000;   
            8'h77: pixels = 12'b000111000000;    
            8'h78: pixels = 12'b001110000000;       
            8'h79: pixels = 12'b001110000000;       
            8'h7A: pixels = 12'b001110000000;     
            8'h7B: pixels = 12'b001110000000;      
            8'h7C: pixels = 12'b001110000000;     
            8'h7D: pixels = 12'b000000000000;         
            8'h7E: pixels = 12'b000000000000;           
            8'h7F: pixels = 12'b000000000000;
            //---------------- ���� 8 -----------------
            8'h80: pixels = 12'b000111111000; 
            8'h81: pixels = 12'b001111111100; 
            8'h82: pixels = 12'b011100011110; 
            8'h83: pixels = 12'b011000001110;
            8'h84: pixels = 12'b011100011110; 
            8'h85: pixels = 12'b001111111100; 
            8'h86: pixels = 12'b001111111100;
            8'h87: pixels = 12'b011100011110; 
            8'h88: pixels = 12'b011000001110; 
            8'h89: pixels = 12'b011000001110; 
            8'h8A: pixels = 12'b011100011110; 
            8'h8B: pixels = 12'b001111111100; 
            8'h8C: pixels = 12'b000111111000; 
            8'h8D: pixels = 12'b000000000000;         
            8'h8E: pixels = 12'b000000000000;        
            8'h8F: pixels = 12'b000000000000; 

            //---------------- ���� 9 -----------------
            8'h90: pixels = 12'b000111111000;  
            8'h91: pixels = 12'b001111111100; 
            8'h92: pixels = 12'b011100011110; 
            8'h93: pixels = 12'b011000001110; 
            8'h94: pixels = 12'b011000001110; 
            8'h95: pixels = 12'b011100011110; 
            8'h96: pixels = 12'b001111111110; 
            8'h97: pixels = 12'b000111111110; 
            8'h98: pixels = 12'b000000001110; 
            8'h99: pixels = 12'b000000001110;
            8'h9A: pixels = 12'b011000011110; 
            8'h9B: pixels = 12'b011111111100; 
            8'h9C: pixels = 12'b001111111000; 
            8'h9D: pixels = 12'b000000000000;            
            8'h9E: pixels = 12'b000000000000;        
            8'h9F: pixels = 12'b000000000000; 

            default: pixels = 12'h000;
        endcase
    end
endmodule